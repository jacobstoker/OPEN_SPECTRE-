remove~!!!
