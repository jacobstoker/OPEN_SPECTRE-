
--   ____  _____  ______ _   _         _____ _____  ______ _____ _______ _____  ______ 
--  / __ \|  __ \|  ____| \ | |       / ____|  __ \|  ____/ ____|__   __|  __ \|  ____|
-- | |  | | |__) | |__  |  \| |      | (___ | |__) | |__ | |       | |  | |__) | |__   
-- | |  | |  ___/|  __| | . ` |       \___ \|  ___/|  __|| |       | |  |  _  /|  __|  
-- | |__| | |    | |____| |\  |       ____) | |    | |___| |____   | |  | | \ \| |____ 
--  \____/|_|    |______|_| \_|      |_____/|_|    |______\_____|  |_|  |_|  \_\______|
--                               ______                                                
--                              |______|                                               
-- Module Name: window_comparator by RD Jordan
-- Created: Early 2023
-- Description: 
-- Dependencies: 
-- Additional Comments: You can view the project here: https://github.com/cfoge/OPEN_SPECTRE-
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity window_comparator is
    Port ( input : in  STD_LOGIC_VECTOR(7 downto 0);
           lower : in  STD_LOGIC_VECTOR(7 downto 0);
           upper : in  STD_LOGIC_VECTOR(7 downto 0);
           output : out  STD_LOGIC);
end window_comparator;

architecture Behavioral of window_comparator is
begin
  output <= '0' when (input < lower) or (input > upper) else '1';
end Behavioral;
