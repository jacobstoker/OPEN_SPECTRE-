package oscillator_pkg is
    constant OSC_PHASE_ACCUMULATOR_WIDTH : integer := 29;
    constant OSC_INDEX_WIDTH             : integer := 10;
    constant OSC_FREQ_CONTROL_WORD_WIDTH : integer := 20;
    constant OSC_AMPLITUDE_WIDTH         : integer := 10;
end package oscillator_pkg;